

module baudRate(clk, outBaud, rst);

    //Define inputs here: 
    input clk; 
    input rst; 

    //Defind outputs here: 
    output reg outBaud; 

    //We know that our internal clock is 100MHz and baudRate is 9600 so we won't try and make this module universal so we can do all math in hosue
    //100M/9600 = 

endmodule